------------------------------------------------------------
-- VHDL CU
-- 2016 9 7 21 24 12
-- Created By "DXP VHDL Generator"
-- "Copyright (c) 2002-2014 Altium Limited"
-- Product Version: 16.1.12.290
------------------------------------------------------------

------------------------------------------------------------
-- VHDL CU
------------------------------------------------------------

Library IEEE;
Use     IEEE.std_logic_1164.all;

Entity CU Is
  port
  (
    CNT_EN : InOut STD_LOGIC;                                -- ObjectKind=Port|PrimaryId=CNT_EN
    CNT_LD : InOut STD_LOGIC;                                -- ObjectKind=Port|PrimaryId=CNT_LD
    DONE   : InOut STD_LOGIC;                                -- ObjectKind=Port|PrimaryId=DONE
    FINI   : InOut STD_LOGIC;                                -- ObjectKind=Port|PrimaryId=FINI
    GO     : InOut STD_LOGIC;                                -- ObjectKind=Port|PrimaryId=GO
    MUX    : InOut STD_LOGIC;                                -- ObjectKind=Port|PrimaryId=MUX
    REG_LD : InOut STD_LOGIC                                 -- ObjectKind=Port|PrimaryId=REG_LD
  );
  attribute MacroCell : boolean;

End CU;
------------------------------------------------------------

------------------------------------------------------------
Architecture Structure Of CU Is


Begin
End Structure;
------------------------------------------------------------

