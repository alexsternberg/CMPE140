////////////////////////////////////////////////////////////////////////////////
// SubModule CMP(GT)
// Created   9/7/2016 10:23:30 PM
////////////////////////////////////////////////////////////////////////////////

module CMP #(parameter width = 32)(B, A, GT);

input [width-1:0] B;
input [width-1:0] A;
output GT;

assign GT = A > B;

endmodule
////////////////////////////////////////////////////////////////////////////////


