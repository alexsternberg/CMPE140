////////////////////////////////////////////////////////////////////////////////
// SubModule BUF
// Created   9/7/2016 10:22:08 PM
////////////////////////////////////////////////////////////////////////////////

module buffer #(parameter width = 32)(
input  [width-1:0] i,
input  oe,
output [width-1:0] o
);

assign o = oe ? i : 'bZ;

endmodule
////////////////////////////////////////////////////////////////////////////////
