////////////////////////////////////////////////////////////////////////////////
// SubModule BUF
// Created   9/7/2016 10:22:08 PM
////////////////////////////////////////////////////////////////////////////////

module BUFFER #(parameter width = 32)(OE, O, I);

input  OE;
output [width-1:0] O;
input  [31:0] I;

assign O = OE ? I : 'bZ;

endmodule
////////////////////////////////////////////////////////////////////////////////
