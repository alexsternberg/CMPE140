////////////////////////////////////////////////////////////////////////////////
// SubModule MUL
// Created   9/7/2016 10:38:20 PM
////////////////////////////////////////////////////////////////////////////////

module MUL #(parameter width = 32)(Z, Y, X);

output [width-1:0] Z;
input  [width-1:0] Y;
input  [width-1:0] X;

assign Z = X * Y;

endmodule
////////////////////////////////////////////////////////////////////////////////
