////////////////////////////////////////////////////////////////////////////////
// SubModule MUX
// Created   9/7/2016 10:33:15 PM
////////////////////////////////////////////////////////////////////////////////

module MUX #(parameter width = 32)(SEL, IN0, IN1, OUT);

input  SEL;
input  [width-1:0] IN0;
input  [width-1:0] IN1;
output [width-1:0] OUT;

assign OUT = SEL ? IN1 : IN0;

endmodule
////////////////////////////////////////////////////////////////////////////////
