////////////////////////////////////////////////////////////////////////////////
// SubModule REGISTER
// Created   9/7/2016 10:25:15 PM
////////////////////////////////////////////////////////////////////////////////

module REGISTER #(parameter width = 32)(LD, CLK, Q, D);

input LD;
input CLK;
input [width-1:0] D;
output [width-1:0] Q;

reg [width-1:0] data;

always@(posedge CLK)
begin
     if(LD) data = D;
end

assign Q = data;

endmodule
////////////////////////////////////////////////////////////////////////////////
