module multiplier(
	input	[31:0] a, b,
	output	[63:0] y);
	
	assign y = a * b;
endmodule
